class yapp_tx_monitor extends uvm_monitor;

  yapp_packet pkt;
  int num_pkt_col;
  virtual interface yapp_if vif;

  uvm_analysis_port #(yapp_packet) item_collected_port;


  `uvm_component_utils_begin(yapp_tx_monitor)
    `uvm_field_int(num_pkt_col, UVM_ALL_ON)
  `uvm_component_utils_end
 
  covergroup yapp_tx_cg with function sample(yapp_packet p);
    option.per_instance = 1; 

    cp_len : coverpoint p.length {
      //bins MIN = {1};
      bins SMALL = {[2:10]};
      bins MEDIUM = {[11:40]};
      bins LARGE = {[41:62]};
      //bins MAX = {63};
    }

    cp_addr : coverpoint p.addr {
      bins LEGAL = {0,1,2};
      //bins ILLEGAL = {3};
      bins ADDR0 = {0};
      bins ADDR1 = {1};
      bins ADDR2 = {2};
    }

    cp_parity_err : coverpoint p.parity_type {
      bins OK  = {GOOD_PARITY};
      bins ERR = {BAD_PARITY};
    }

    cross_len_addr_par : cross cp_len, cp_addr, cp_parity_err {
      //ignore_bins illegal_addr = binsof(cp_addr.ILLEGAL);
      //ignore_bins ok_parity    = binsof(cp_parity_err.OK);
    }

  endgroup

  function new (string name , uvm_component parent);
    super.new(name, parent);
    item_collected_port = new("item_collected_port", this);
    yapp_tx_cg = new();
  endfunction: new

  function void connect_phase(uvm_phase phase);
    if (!yapp_vif_config::get(this, get_full_name(),"vif",vif))
      `uvm_error("NOVIF", {"Virtual interface must be set for:", get_full_name(), " .vif"})
  endfunction:connect_phase

  // UVM run() phase
  task run_phase(uvm_phase phase);
    // Look for packets after reset
    @(posedge vif.reset)
    @(negedge vif.reset)
    `uvm_info(get_type_name(), "Detected Reset Done", UVM_MEDIUM)
    forever begin 
      // Create collected packet instance
      pkt = yapp_packet::type_id::create("pkt", this);

      // concurrent blocks for packet collection and transaction recording
      fork
        // collect packet
        vif.collect_packet(pkt.length, pkt.addr, pkt.payload, pkt.parity);
        // trigger transaction at start of packet
        @(posedge vif.monstart) void'(begin_tr(pkt, "Monitor_YAPP_Packet"));
      join

      pkt.parity_type = (pkt.parity == pkt.calc_parity()) ? GOOD_PARITY : BAD_PARITY;


      yapp_tx_cg.sample(pkt);
      end_tr(pkt);

      `uvm_info(get_type_name(), $sformatf("Packet Collected :\n%s", pkt.sprint()), UVM_LOW)
      item_collected_port.write(pkt);
      num_pkt_col++;
    end
  endtask : run_phase





  // UVM report_phase
  function void report_phase(uvm_phase phase);
    `uvm_info(get_type_name(), $sformatf("Report: YAPP Monitor Collected %0d Packets", num_pkt_col), UVM_LOW)
  endfunction : report_phase

endclass: yapp_tx_monitor
